`timescale 1ns/1ps

`include "../../lib/std/std_util.svh"
`include "../../lib/std/std_mem.svh"

`include "../../lib/isa/rv.svh"
`include "../../lib/isa/rv32.svh"
`include "../../lib/isa/rv32i.svh"

`include "../../lib/gecko/gecko.svh"

module gecko_micro_tb
    import rv::*;
    import rv32::*;
    import rv32i::*;
    import gecko::*;
#()();

    logic clk, rst;
    clk_rst_gen clk_rst_gen_inst(.clk, .rst);

    logic faulted_flag, finished_flag;

    gecko_micro #(
        .INST_LATENCY(1),
        .DATA_LATENCY(1)
    ) gecko_micro_inst (
        .clk, .rst,
        .faulted_flag, .finished_flag
    );

endmodule
