`ifndef __AXI4_STREAM__
`define __AXI4_STREAM__

package axi4_stream;

endpackage

`endif
