`timescale 1ns/1ps

`ifdef __LINTER__

`include "../../lib/std/std_util.svh"
`include "../../lib/isa/rv.svh"
`include "../../lib/isa/rv32.svh"
`include "../../lib/isa/rv32f.svh"
`include "../../lib/fpu/fpu.svh"
`include "../../lib/fpu/fpu_add.svh"
`include "../../lib/basilisk/basilisk.svh"

`else

`include "std_util.svh"
`include "rv.svh"
`include "rv32.svh"
`include "rv32f.svh"
`include "basilisk.svh"
`include "fpu.svh"
`include "fpu_add.svh"

`endif

module basilisk_add_exponent
    import rv::*;
    import rv32::*;
    import rv32f::*;
    import fpu::*;
    import fpu_add::*;
    import basilisk::*;
#(
    parameter int OUTPUT_REGISTER_MODE = 1
)(
    input logic clk, rst,

    std_stream_intf.in add_command, // basilisk_add_command_t
    std_stream_intf.in mult_add_command, // basilisk_add_command_t
    std_stream_intf.out add_exponent_command // fpu_add_exp_result_t
);

    std_stream_intf #(.T(fpu_add_exp_result_t)) next_add_exponent_command (.clk, .rst);

    logic enable, consume_add, consume_mult_add, produce;

    std_flow_lite #(
        .NUM_INPUTS(2),
        .NUM_OUTPUTS(1)
    ) std_flow_lite_inst (
        .clk, .rst,

        .valid_input({add_command.valid, mult_add_command.valid}),
        .ready_input({add_command.ready, mult_add_command.ready}),

        .valid_output({next_add_exponent_command.valid}),
        .ready_output({next_add_exponent_command.ready}),

        .consume({consume_add, consume_mult_add}),
        .produce,
        .enable
    );

    std_flow_stage #(
        .T(fpu_add_exp_result_t),
        .MODE(OUTPUT_REGISTER_MODE)
    ) output_stage_inst (
        .clk, .rst,
        .stream_in(next_add_exponent_command), .stream_out(add_exponent_command)
    );

    always_comb begin
        automatic basilisk_add_command_t chosen_command;

        consume_add = 'b1;
        consume_mult_add = 'b0;
        produce = 'b1;

        if (mult_add_command.valid) begin
            consume_mult_add = 'b1;
            consume_add = 'b0;
            chosen_command = basilisk_add_command_t'(mult_add_command.payload);
        end else begin
            chosen_command = basilisk_add_command_t'(add_command.payload);
        end

        next_add_exponent_command.payload = fpu_float_add_exponent(
                chosen_command.a, chosen_command.b,
                chosen_command.conditions_a, chosen_command.conditions_b,
                chosen_command.mode
        );
    end

endmodule
