`ifndef __RV_AXI4_DEF__
`define __RV_AXI4_DEF__

/*
 * Write Address Defines
 */

`define RV_AXI4_AW_PORTS_OUT(PREFIX, ADDR_WIDTH, DATA_WIDTH, ID_WIDTH, USER_WIDTH) \
    `RV_AXI4_AW_PORTS(output, input, PREFIX, ADDR_WIDTH, DATA_WIDTH, ID_WIDTH, USER_WIDTH)
`define RV_AXI4_AW_PORTS_IN(PREFIX, ADDR_WIDTH, DATA_WIDTH, ID_WIDTH, USER_WIDTH) \
    `RV_AXI4_AW_PORTS(input, output, PREFIX, ADDR_WIDTH, DATA_WIDTH, ID_WIDTH, USER_WIDTH)
`define RV_AXI4_AW_PORTS(FLOW_DIR, BACKFLOW_DIR, PREFIX, ADDR_WIDTH, DATA_WIDTH, ID_WIDTH, USER_WIDTH) \
    FLOW_DIR wire ``PREFIX``_AWVALID, BACKFLOW_DIR wire ``PREFIX``_AWREADY, \
    FLOW_DIR wire [ADDR_WIDTH-1:0] ``PREFIX``_AWADDR, \
    FLOW_DIR wire [1:0]            ``PREFIX``_AWBURST, \
    FLOW_DIR wire [3:0]            ``PREFIX``_AWCACHE, \
    FLOW_DIR wire [7:0]            ``PREFIX``_AWLEN, \
    FLOW_DIR wire                  ``PREFIX``_AWLOCK, \
    FLOW_DIR wire [2:0]            ``PREFIX``_AWPROT, \
    FLOW_DIR wire [3:0]            ``PREFIX``_AWQOS, \
    FLOW_DIR wire [2:0]            ``PREFIX``_AWSIZE, \
    FLOW_DIR wire [USER_WIDTH-1:0] ``PREFIX``_AWUSER, \
    FLOW_DIR wire [ID_WIDTH-1:0]   ``PREFIX``_AWID

`define RV_AXI4_AW_CONNECT(PREFIX_IN, PREFIX_OUT) \
    assign ``PREFIX_OUT``AWVALID = ``PREFIX_IN``AWVALID; \
    assign ``PREFIX_IN``AWREADY  = ``PREFIX_OUT``AWREADY; \
    assign ``PREFIX_OUT``AWADDR  = ``PREFIX_IN``AWADDR; \
    assign ``PREFIX_OUT``AWBURST = rv_axi4::rv_axi4_burst'(``PREFIX_IN``AWBURST); \
    assign ``PREFIX_OUT``AWCACHE = rv_axi4::rv_axi4_cache'(``PREFIX_IN``AWCACHE); \
    assign ``PREFIX_OUT``AWLEN   = ``PREFIX_IN``AWLEN; \
    assign ``PREFIX_OUT``AWLOCK  = rv_axi4::rv_axi4_lock'(``PREFIX_IN``AWLOCK); \
    assign ``PREFIX_OUT``AWPROT  = rv_axi4::rv_axi4_prot'(``PREFIX_IN``AWPROT); \
    assign ``PREFIX_OUT``AWQOS   = ``PREFIX_IN``AWQOS; \
    assign ``PREFIX_OUT``AWSIZE  = ``PREFIX_IN``AWSIZE; \
    assign ``PREFIX_OUT``AWUSER  = ``PREFIX_IN``AWUSER; \
    assign ``PREFIX_OUT``AWID    = ``PREFIX_IN``AWID;

`define RV_AXI4_AW_CONNECT_PORTS(PREFIX_IN, PREFIX_OUT) \
    .``PREFIX_OUT``AWVALID(``PREFIX_IN``AWVALID), \
    .``PREFIX_OUT``AWREADY(``PREFIX_IN``AWREADY), \
    .``PREFIX_OUT``AWADDR(``PREFIX_IN``AWADDR), \
    .``PREFIX_OUT``AWBURST(``PREFIX_IN``AWBURST), \
    .``PREFIX_OUT``AWCACHE(``PREFIX_IN``AWCACHE), \
    .``PREFIX_OUT``AWLEN(``PREFIX_IN``AWLEN), \
    .``PREFIX_OUT``AWLOCK(``PREFIX_IN``AWLOCK), \
    .``PREFIX_OUT``AWPROT(``PREFIX_IN``AWPROT), \
    .``PREFIX_OUT``AWQOS(``PREFIX_IN``AWQOS), \
    .``PREFIX_OUT``AWSIZE(``PREFIX_IN``AWSIZE), \
    .``PREFIX_OUT``AWUSER(``PREFIX_IN``AWUSER), \
    .``PREFIX_OUT``AWID(``PREFIX_IN``AWID)

/*
 * Write Data Defines
 */

`define RV_AXI4_W_PORTS_OUT(PREFIX, ADDR_WIDTH, DATA_WIDTH, ID_WIDTH, USER_WIDTH) \
    `RV_AXI4_W_PORTS(output, input, PREFIX, ADDR_WIDTH, DATA_WIDTH, ID_WIDTH, USER_WIDTH)
`define RV_AXI4_W_PORTS_IN(PREFIX, ADDR_WIDTH, DATA_WIDTH, ID_WIDTH, USER_WIDTH) \
    `RV_AXI4_W_PORTS(input, output, PREFIX, ADDR_WIDTH, DATA_WIDTH, ID_WIDTH, USER_WIDTH)
`define RV_AXI4_W_PORTS(FLOW_DIR, BACKFLOW_DIR, PREFIX, ADDR_WIDTH, DATA_WIDTH, ID_WIDTH, USER_WIDTH) \
    FLOW_DIR wire ``PREFIX``_WVALID, BACKFLOW_DIR wire ``PREFIX``_WREADY, \
    FLOW_DIR wire [DATA_WIDTH-1:0]     ``PREFIX``_WDATA, \
    FLOW_DIR wire [(DATA_WIDTH/8)-1:0] ``PREFIX``_WSTRB, \
    FLOW_DIR wire                      ``PREFIX``_WLAST

`define RV_AXI4_W_CONNECT(PREFIX_IN, PREFIX_OUT) \
    assign ``PREFIX_OUT``WVALID = ``PREFIX_IN``WVALID; \
    assign ``PREFIX_IN``WREADY  = ``PREFIX_OUT``WREADY; \
    assign ``PREFIX_OUT``WDATA  = ``PREFIX_IN``WDATA; \
    assign ``PREFIX_OUT``WSTRB  = ``PREFIX_IN``WSTRB; \
    assign ``PREFIX_OUT``WLAST  = ``PREFIX_IN``WLAST;

`define RV_AXI4_W_CONNECT_PORTS(PREFIX_IN, PREFIX_OUT) \
    .``PREFIX_OUT``WVALID(``PREFIX_IN``WVALID), \
    .``PREFIX_OUT``WREADY(``PREFIX_IN``WREADY), \
    .``PREFIX_OUT``WDATA(``PREFIX_IN``WDATA), \
    .``PREFIX_OUT``WSTRB(``PREFIX_IN``WSTRB), \
    .``PREFIX_OUT``WLAST(``PREFIX_IN``WLAST)

/*
 * Write Respond Defines
 */

`define RV_AXI4_B_PORTS_OUT(PREFIX, ADDR_WIDTH, DATA_WIDTH, ID_WIDTH, USER_WIDTH) \
    `RV_AXI4_B_PORTS(output, input, PREFIX, ADDR_WIDTH, DATA_WIDTH, ID_WIDTH, USER_WIDTH)
`define RV_AXI4_B_PORTS_IN(PREFIX, ADDR_WIDTH, DATA_WIDTH, ID_WIDTH, USER_WIDTH) \
    `RV_AXI4_B_PORTS(input, output, PREFIX, ADDR_WIDTH, DATA_WIDTH, ID_WIDTH, USER_WIDTH)
`define RV_AXI4_B_PORTS(FLOW_DIR, BACKFLOW_DIR, PREFIX, ADDR_WIDTH, DATA_WIDTH, ID_WIDTH, USER_WIDTH) \
    FLOW_DIR wire ``PREFIX``_BVALID, BACKFLOW_DIR wire ``PREFIX``_BREADY, \
    FLOW_DIR wire [1:0]          ``PREFIX``_BRESP, \
    FLOW_DIR wire [ID_WIDTH-1:0] ``PREFIX``_BID

`define RV_AXI4_B_CONNECT(PREFIX_IN, PREFIX_OUT) \
    assign ``PREFIX_OUT``BVALID = ``PREFIX_IN``BVALID; \
    assign ``PREFIX_IN``BREADY  = ``PREFIX_OUT``BREADY; \
    assign ``PREFIX_OUT``BRESP  = rv_axi4::rv_axi4_resp'(``PREFIX_IN``BRESP); \
    assign ``PREFIX_OUT``BID    = ``PREFIX_IN``BID;

`define RV_AXI4_B_CONNECT_PORTS(PREFIX_IN, PREFIX_OUT) \
    .``PREFIX_OUT``BVALID(``PREFIX_IN``BVALID), \
    .``PREFIX_OUT``BREADY(``PREFIX_IN``BREADY), \
    .``PREFIX_OUT``BRESP(``PREFIX_IN``BRESP), \
    .``PREFIX_OUT``BID(``PREFIX_IN``BID)

/*
 * Read Address Defines
 */

`define RV_AXI4_AR_PORTS_OUT(PREFIX, ADDR_WIDTH, DATA_WIDTH, ID_WIDTH, USER_WIDTH) \
    `RV_AXI4_AR_PORTS(output, input, PREFIX, ADDR_WIDTH, DATA_WIDTH, ID_WIDTH, USER_WIDTH)
`define RV_AXI4_AR_PORTS_IN(PREFIX, ADDR_WIDTH, DATA_WIDTH, ID_WIDTH, USER_WIDTH) \
    `RV_AXI4_AR_PORTS(input, output, PREFIX, ADDR_WIDTH, DATA_WIDTH, ID_WIDTH, USER_WIDTH)
`define RV_AXI4_AR_PORTS(FLOW_DIR, BACKFLOW_DIR, PREFIX, ADDR_WIDTH, DATA_WIDTH, ID_WIDTH, USER_WIDTH) \
    FLOW_DIR wire ``PREFIX``_ARVALID, BACKFLOW_DIR wire ``PREFIX``_ARREADY, \
    FLOW_DIR wire [ADDR_WIDTH-1:0] ``PREFIX``_ARADDR, \
    FLOW_DIR wire [1:0]            ``PREFIX``_ARBURST, \
    FLOW_DIR wire [3:0]            ``PREFIX``_ARCACHE, \
    FLOW_DIR wire [7:0]            ``PREFIX``_ARLEN, \
    FLOW_DIR wire                  ``PREFIX``_ARLOCK, \
    FLOW_DIR wire [2:0]            ``PREFIX``_ARPROT, \
    FLOW_DIR wire [3:0]            ``PREFIX``_ARQOS, \
    FLOW_DIR wire [2:0]            ``PREFIX``_ARSIZE, \
    FLOW_DIR wire [USER_WIDTH-1:0] ``PREFIX``_ARUSER, \
    FLOW_DIR wire [ID_WIDTH-1:0]   ``PREFIX``_ARID

`define RV_AXI4_AR_CONNECT(PREFIX_IN, PREFIX_OUT) \
    assign ``PREFIX_OUT``ARVALID = ``PREFIX_IN``ARVALID; \
    assign ``PREFIX_IN``ARREADY  = ``PREFIX_OUT``ARREADY; \
    assign ``PREFIX_OUT``ARADDR  = ``PREFIX_IN``ARADDR; \
    assign ``PREFIX_OUT``ARBURST = rv_axi4::rv_axi4_burst'(``PREFIX_IN``ARBURST); \
    assign ``PREFIX_OUT``ARCACHE = rv_axi4::rv_axi4_cache'(``PREFIX_IN``ARCACHE); \
    assign ``PREFIX_OUT``ARLEN   = ``PREFIX_IN``ARLEN; \
    assign ``PREFIX_OUT``ARLOCK  = rv_axi4::rv_axi4_lock'(``PREFIX_IN``ARLOCK); \
    assign ``PREFIX_OUT``ARPROT  = rv_axi4::rv_axi4_prot'(``PREFIX_IN``ARPROT); \
    assign ``PREFIX_OUT``ARQOS   = ``PREFIX_IN``ARQOS; \
    assign ``PREFIX_OUT``ARSIZE  = ``PREFIX_IN``ARSIZE; \
    assign ``PREFIX_OUT``ARUSER  = ``PREFIX_IN``ARUSER; \
    assign ``PREFIX_OUT``ARID    = ``PREFIX_IN``ARID;

`define RV_AXI4_AR_CONNECT_PORTS(PREFIX_IN, PREFIX_OUT) \
    .``PREFIX_OUT``ARVALID(``PREFIX_IN``ARVALID), \
    .``PREFIX_OUT``ARREADY(``PREFIX_IN``ARREADY), \
    .``PREFIX_OUT``ARADDR(``PREFIX_IN``ARADDR), \
    .``PREFIX_OUT``ARBURST(``PREFIX_IN``ARBURST), \
    .``PREFIX_OUT``ARCACHE(``PREFIX_IN``ARCACHE), \
    .``PREFIX_OUT``ARLEN(``PREFIX_IN``ARLEN), \
    .``PREFIX_OUT``ARLOCK(``PREFIX_IN``ARLOCK), \
    .``PREFIX_OUT``ARPROT(``PREFIX_IN``ARPROT), \
    .``PREFIX_OUT``ARQOS(``PREFIX_IN``ARQOS), \
    .``PREFIX_OUT``ARSIZE(``PREFIX_IN``ARSIZE), \
    .``PREFIX_OUT``ARUSER(``PREFIX_IN``ARUSER), \
    .``PREFIX_OUT``ARID(``PREFIX_IN``ARID)

/*
 * Read Data Defines
 */

`define RV_AXI4_R_PORTS_OUT(PREFIX, ADDR_WIDTH, DATA_WIDTH, ID_WIDTH, USER_WIDTH) \
    `RV_AXI4_R_PORTS(output, input, PREFIX, ADDR_WIDTH, DATA_WIDTH, ID_WIDTH, USER_WIDTH)
`define RV_AXI4_R_PORTS_IN(PREFIX, ADDR_WIDTH, DATA_WIDTH, ID_WIDTH, USER_WIDTH) \
    `RV_AXI4_R_PORTS(input, output, PREFIX, ADDR_WIDTH, DATA_WIDTH, ID_WIDTH, USER_WIDTH)
`define RV_AXI4_R_PORTS(FLOW_DIR, BACKFLOW_DIR, PREFIX, ADDR_WIDTH, DATA_WIDTH, ID_WIDTH, USER_WIDTH) \
    FLOW_DIR wire ``PREFIX``_RVALID, BACKFLOW_DIR wire ``PREFIX``_RREADY, \
    FLOW_DIR wire [DATA_WIDTH-1:0] ``PREFIX``_RDATA, \
    FLOW_DIR wire                  ``PREFIX``_RLAST, \
    FLOW_DIR wire [1:0]            ``PREFIX``_RRESP, \
    FLOW_DIR wire [ID_WIDTH-1:0]   ``PREFIX``_RID

`define RV_AXI4_R_CONNECT(PREFIX_IN, PREFIX_OUT) \
    assign ``PREFIX_OUT``RVALID = ``PREFIX_IN``RVALID; \
    assign ``PREFIX_IN``RREADY  = ``PREFIX_OUT``RREADY; \
    assign ``PREFIX_OUT``RDATA  = ``PREFIX_IN``RDATA; \
    assign ``PREFIX_OUT``RLAST  = ``PREFIX_IN``RLAST; \
    assign ``PREFIX_OUT``RRESP  = rv_axi4::rv_axi4_resp'(``PREFIX_IN``RRESP); \
    assign ``PREFIX_OUT``RID    = ``PREFIX_IN``RID;

`define RV_AXI4_R_CONNECT_PORTS(PREFIX_IN, PREFIX_OUT) \
    .``PREFIX_OUT``RVALID(``PREFIX_IN``RVALID), \
    .``PREFIX_OUT``RREADY(``PREFIX_IN``RREADY), \
    .``PREFIX_OUT``RDATA(``PREFIX_IN``RDATA), \
    .``PREFIX_OUT``RLAST(``PREFIX_IN``RLAST), \
    .``PREFIX_OUT``RRESP(``PREFIX_IN``RRESP), \
    .``PREFIX_OUT``RID(``PREFIX_IN``RID)

/*
 * Entire AXI4 Bus Definitions
 */

`define RV_AXI4_PORTS_MASTER(PREFIX, ADDR_WIDTH, DATA_WIDTH, ID_WIDTH, USER_WIDTH) \
    `RV_AXI4_AW_PORTS_OUT(PREFIX, ADDR_WIDTH, DATA_WIDTH, ID_WIDTH, USER_WIDTH), \
    `RV_AXI4_W_PORTS_OUT(PREFIX, ADDR_WIDTH, DATA_WIDTH, ID_WIDTH, USER_WIDTH), \
    `RV_AXI4_B_PORTS_IN(PREFIX, ADDR_WIDTH, DATA_WIDTH, ID_WIDTH, USER_WIDTH), \
    `RV_AXI4_AR_PORTS_OUT(PREFIX, ADDR_WIDTH, DATA_WIDTH, ID_WIDTH, USER_WIDTH), \
    `RV_AXI4_R_PORTS_IN(PREFIX, ADDR_WIDTH, DATA_WIDTH, ID_WIDTH, USER_WIDTH)

`define RV_AXI4_PORTS_SLAVE(PREFIX, ADDR_WIDTH, DATA_WIDTH, ID_WIDTH, USER_WIDTH) \
    `RV_AXI4_AW_PORTS_IN(PREFIX, ADDR_WIDTH, DATA_WIDTH, ID_WIDTH, USER_WIDTH), \
    `RV_AXI4_W_PORTS_IN(PREFIX, ADDR_WIDTH, DATA_WIDTH, ID_WIDTH, USER_WIDTH), \
    `RV_AXI4_B_PORTS_OUT(PREFIX, ADDR_WIDTH, DATA_WIDTH, ID_WIDTH, USER_WIDTH), \
    `RV_AXI4_AR_PORTS_IN(PREFIX, ADDR_WIDTH, DATA_WIDTH, ID_WIDTH, USER_WIDTH), \
    `RV_AXI4_R_PORTS_OUT(PREFIX, ADDR_WIDTH, DATA_WIDTH, ID_WIDTH, USER_WIDTH)

`define RV_AXI4_INTF_MASTER(PREFIX) \
    rv_axi4_aw_intf.out ``PREFIX``_aw, \
    rv_axi4_w_intf.out ``PREFIX``_w, \
    rv_axi4_b_intf.in ``PREFIX``_b, \
    rv_axi4_ar_intf.out ``PREFIX``_ar, \
    rv_axi4_r_intf.in ``PREFIX``_r

`define RV_AXI4_INTF_SLAVE(PREFIX) \
    rv_axi4_aw_intf.in ``PREFIX``_aw, \
    rv_axi4_w_intf.in ``PREFIX``_w, \
    rv_axi4_b_intf.out ``PREFIX``_b, \
    rv_axi4_ar_intf.in ``PREFIX``_ar, \
    rv_axi4_r_intf.out ``PREFIX``_r

`define RV_AXI4_CREATE_INTF(PREFIX, AW, DW, IW, UW) \
    rv_axi4_aw_intf #(.ADDR_WIDTH(AW), .USER_WIDTH(UW), .ID_WIDTH(IW)) ``PREFIX``_aw (); \
    rv_axi4_w_intf #(.DATA_WIDTH(DW))                                  ``PREFIX``_w (); \
    rv_axi4_b_intf #(.ID_WIDTH(IW))                                    ``PREFIX``_b (); \
    rv_axi4_ar_intf #(.ADDR_WIDTH(AW), .USER_WIDTH(UW), .ID_WIDTH(IW)) ``PREFIX``_ar (); \
    rv_axi4_r_intf #(.DATA_WIDTH(DW), .ID_WIDTH(IW))                   ``PREFIX``_r ();

`define RV_AXI4_CONNECT(PREFIX_IN, PREFIX_OUT) \
    `RV_AXI4_AW_CONNECT(PREFIX_IN, PREFIX_OUT) \
    `RV_AXI4_W_CONNECT(PREFIX_IN, PREFIX_OUT) \
    `RV_AXI4_B_CONNECT(PREFIX_OUT, PREFIX_IN) \
    `RV_AXI4_AR_CONNECT(PREFIX_IN, PREFIX_OUT) \
    `RV_AXI4_R_CONNECT(PREFIX_OUT, PREFIX_IN)

`define RV_AXI4_CONNECT_PORTS_TO_INTF(PREFIX_IN, PREFIX_OUT) \
    `RV_AXI4_AW_CONNECT(``PREFIX_IN``_, ``PREFIX_OUT``_aw.) \
    `RV_AXI4_W_CONNECT(``PREFIX_IN``_, ``PREFIX_OUT``_w.) \
    `RV_AXI4_B_CONNECT(``PREFIX_OUT``_b., ``PREFIX_IN``_) \
    `RV_AXI4_AR_CONNECT(``PREFIX_IN``_, ``PREFIX_OUT``_ar.) \
    `RV_AXI4_R_CONNECT(``PREFIX_OUT``_r., ``PREFIX_IN``_)

`define RV_AXI4_CONNECT_INTF_TO_PORTS(PREFIX_IN, PREFIX_OUT) \
    `RV_AXI4_AW_CONNECT(``PREFIX_IN``_aw., ``PREFIX_OUT``_) \
    `RV_AXI4_W_CONNECT(``PREFIX_IN``_w., ``PREFIX_OUT``_) \
    `RV_AXI4_B_CONNECT(``PREFIX_OUT``_, ``PREFIX_IN``_b.) \
    `RV_AXI4_AR_CONNECT(``PREFIX_IN``_ar., ``PREFIX_OUT``_) \
    `RV_AXI4_R_CONNECT(``PREFIX_OUT``_, ``PREFIX_IN``_r.)

`define RV_AXI4_CONNECT_PORTS(PREFIX_IN, PREFIX_OUT) \
    `RV_AXI4_AW_CONNECT_PORTS(``PREFIX_IN``_, ``PREFIX_OUT``_), \
    `RV_AXI4_W_CONNECT_PORTS(``PREFIX_IN``_, ``PREFIX_OUT``_), \
    `RV_AXI4_B_CONNECT_PORTS(``PREFIX_IN``_, ``PREFIX_OUT``_), \
    `RV_AXI4_AR_CONNECT_PORTS(``PREFIX_IN``_, ``PREFIX_OUT``_), \
    `RV_AXI4_R_CONNECT_PORTS(``PREFIX_IN``_, ``PREFIX_OUT``_)

`endif
