package axi4_stream_pkg;

endpackage
