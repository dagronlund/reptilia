`ifndef __RV_CACHE__
`define __RV_CACHE__

package rv_cache;

endpackage

`endif
