`ifndef __RV32F__
`define __RV32F__

`ifdef __SIMULATION__
`include "rv.svh"
`include "rv32.svh"
`endif

package rv32f;

    import rv::*;
    import rv32::*;

endpackage

`endif
