`ifndef __RV32_CSR__
`define __RV32_CSR__

package rv32_csr;

endpackage

`endif
